** Profile: "SCHEMATIC1-NCS2200"  [ C:\ON-Semi\NCS2200\PSPICE\ncs2200-schematic1-ncs2200.sim ] 

** Creating circuit file "ncs2200-schematic1-ncs2200.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB ".\ncs2200p.lib" 
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2ms 0 0.1m 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\ncs2200-SCHEMATIC1.net" 


.END
