** Profile: "SCHEMATIC1-Exam_8_1"  [ D:\Ian_Jung\workplace\PSpice\Exam_8_1-PSpiceFiles\SCHEMATIC1\Exam_8_1.sim ] 

** Creating circuit file "Exam_8_1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 50m 0 
.MC 100 TRAN V(out0 YMAX OUTPUT ALL SEED=43 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
