** Profile: "SCHEMATIC1-BJT_Amp"  [ D:\Ian_Jung\workplace\PSpice\NPN_1-PSpiceFiles\SCHEMATIC1\BJT_Amp.sim ] 

** Creating circuit file "BJT_Amp.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 1 10meg
.NOISE V([OUT]) V_Vsig 10
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
