** Profile: "SCHEMATIC1-IV_curve"  [ D:\Ian_Jung\workplace\PSpice\FET_AMP_2-PSpiceFiles\SCHEMATIC1\IV_curve.sim ] 

** Creating circuit file "IV_curve.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_VDS 0 5 0.01 
+ LIN V_VGS 0 2 0.05 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
