** Profile: "SCHEMATIC1-Tran"  [ D:\Ian_Jung\workplace\PSpice\Timer_555-PSpiceFiles\SCHEMATIC1\Tran.sim ] 

** Creating circuit file "Tran.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../library/ncs2200p.lib" 
.LIB "../../../library/cmos_nor_gate.lib" 
.LIB "../../../library/cmos_inv.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2m 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
