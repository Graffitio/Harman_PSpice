** Profile: "SCHEMATIC1-BJT_IV_cur"  [ D:\Ian_Jung\workplace\PSpice\NPN_IV_cur-PSpiceFiles\SCHEMATIC1\BJT_IV_cur.sim ] 

** Creating circuit file "BJT_IV_cur.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V1 0 5V 0.0005 
.STEP LIN I_I1 0 100u 20u 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
