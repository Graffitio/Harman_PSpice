** Profile: "SCHEMATIC1-Counter"  [ D:\Ian_Jung\workplace\PSpice\Counter-PSpiceFiles\SCHEMATIC1\Counter.sim ] 

** Creating circuit file "Counter.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10us 0 1n 
.OPTIONS ADVCONV
.OPTIONS DIGINITSTATE= 1
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
