** Profile: "SCHEMATIC1-BP_test1"  [ D:\Ian_Jung\workplace\PSpice\part_3_bias_point-PSpiceFiles\SCHEMATIC1\BP_test1.sim ] 

** Creating circuit file "BP_test1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.SENS V([OUT]) 
.TF V(R_R2) V_V1
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
